library verilog;
use verilog.vl_types.all;
entity Celda_vlg_vec_tst is
end Celda_vlg_vec_tst;
