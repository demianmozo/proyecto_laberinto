library verilog;
use verilog.vl_types.all;
entity decido_accion_vlg_vec_tst is
end decido_accion_vlg_vec_tst;
