library verilog;
use verilog.vl_types.all;
entity seleccionadores_mux_vlg_vec_tst is
end seleccionadores_mux_vlg_vec_tst;
