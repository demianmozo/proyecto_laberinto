library verilog;
use verilog.vl_types.all;
entity Matriz_ubicacion_vlg_vec_tst is
end Matriz_ubicacion_vlg_vec_tst;
