library verilog;
use verilog.vl_types.all;
entity SENT_ACTUAL_vlg_vec_tst is
end SENT_ACTUAL_vlg_vec_tst;
