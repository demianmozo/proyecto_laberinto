library verilog;
use verilog.vl_types.all;
entity Control_Motores_vlg_vec_tst is
end Control_Motores_vlg_vec_tst;
