-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Jul 28 00:11:18 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Motores IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SR : IN STD_LOGIC := '0';
        SL : IN STD_LOGIC := '0';
        SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        fin_giro : IN STD_LOGIC := '0';
        llego : IN STD_LOGIC := '0';
        MD0 : OUT STD_LOGIC;
        MI0 : OUT STD_LOGIC;
        MD1 : OUT STD_LOGIC;
        MI1 : OUT STD_LOGIC;
        h_giro : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END Motores;

ARCHITECTURE BEHAVIOR OF Motores IS
    TYPE type_fstate IS (Avanza,Corrige_izq,Corrige_der,Gira_90_izq,Gira_90_der,Gira_180,Ganamos);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= Avanza;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,SR,SL,SEL,fin_giro,llego)
    BEGIN
        MD0 <= '0';
        MI0 <= '0';
        MD1 <= '0';
        MI1 <= '0';
        h_giro <= "00";
        CASE fstate IS
            WHEN Avanza =>
                IF (((((SEL(1 DOWNTO 0) = "00") AND (SR = '1')) AND (SL = '1')) AND (llego = '0'))) THEN
                    reg_fstate <= Avanza;
                ELSIF (((((SEL(1 DOWNTO 0) = "00") AND (SR = '0')) AND (SL = '1')) AND (llego = '0'))) THEN
                    reg_fstate <= Corrige_izq;
                ELSIF (((((SEL(1 DOWNTO 0) = "00") AND (SR = '1')) AND (SL = '0')) AND (llego = '0'))) THEN
                    reg_fstate <= Corrige_der;
                ELSIF (((SEL(1 DOWNTO 0) = "01") AND (llego = '0'))) THEN
                    reg_fstate <= Gira_90_izq;
                ELSIF (((SEL(1 DOWNTO 0) = "10") AND (llego = '0'))) THEN
                    reg_fstate <= Gira_90_der;
                ELSIF (((SEL(1 DOWNTO 0) = "11") AND (llego = '0'))) THEN
                    reg_fstate <= Gira_180;
                ELSIF ((llego = '1')) THEN
                    reg_fstate <= Ganamos;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Avanza;
                END IF;

                MD0 <= '1';

                MI0 <= '1';

                MD1 <= '0';

                h_giro <= "00";

                MI1 <= '0';
            WHEN Corrige_izq =>
                IF ((((SR = '0') AND (SEL(1 DOWNTO 0) = "00")) AND (llego = '0'))) THEN
                    reg_fstate <= Corrige_izq;
                ELSIF ((((SR = '1') AND (SEL(1 DOWNTO 0) = "00")) AND (llego = '0'))) THEN
                    reg_fstate <= Avanza;
                ELSIF ((llego = '1')) THEN
                    reg_fstate <= Ganamos;
                ELSIF ((((SR = '0') AND (SEL(1 DOWNTO 0) = "01")) AND (llego = '0'))) THEN
                    reg_fstate <= Gira_90_izq;
                ELSIF ((((SR = '0') AND (SEL(1 DOWNTO 0) = "10")) AND (llego = '0'))) THEN
                    reg_fstate <= Gira_90_der;
                ELSIF ((((SR = '0') AND (SEL(1 DOWNTO 0) = "11")) AND (llego = '0'))) THEN
                    reg_fstate <= Gira_180;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Corrige_izq;
                END IF;

                MD0 <= '1';

                MI0 <= '0';

                MD1 <= '0';

                h_giro <= "00";

                MI1 <= '0';
            WHEN Corrige_der =>
                IF ((((SL = '0') AND (SEL(1 DOWNTO 0) = "00")) AND (llego = '0'))) THEN
                    reg_fstate <= Corrige_der;
                ELSIF ((((SL = '1') AND (SEL(1 DOWNTO 0) = "00")) AND (llego = '0'))) THEN
                    reg_fstate <= Avanza;
                ELSIF ((llego = '1')) THEN
                    reg_fstate <= Ganamos;
                ELSIF ((((SL = '0') AND (SEL(1 DOWNTO 0) = "01")) AND (llego = '0'))) THEN
                    reg_fstate <= Gira_90_izq;
                ELSIF ((((SL = '0') AND (SEL(1 DOWNTO 0) = "10")) AND (llego = '0'))) THEN
                    reg_fstate <= Gira_90_der;
                ELSIF ((((SL = '0') AND (SEL(1 DOWNTO 0) = "11")) AND (llego = '0'))) THEN
                    reg_fstate <= Gira_180;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Corrige_der;
                END IF;

                MD0 <= '0';

                MI0 <= '1';

                MD1 <= '0';

                h_giro <= "00";

                MI1 <= '0';
            WHEN Gira_90_izq =>
                IF ((fin_giro = '0')) THEN
                    reg_fstate <= Gira_90_izq;
                ELSIF ((fin_giro = '1')) THEN
                    reg_fstate <= Avanza;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Gira_90_izq;
                END IF;

                MD0 <= '1';

                MI0 <= '0';

                MD1 <= '0';

                h_giro <= "01";

                MI1 <= '1';
            WHEN Gira_90_der =>
                IF ((fin_giro = '0')) THEN
                    reg_fstate <= Gira_90_der;
                ELSIF ((fin_giro = '1')) THEN
                    reg_fstate <= Avanza;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Gira_90_der;
                END IF;

                MD0 <= '0';

                MI0 <= '1';

                MD1 <= '1';

                h_giro <= "01";

                MI1 <= '0';
            WHEN Gira_180 =>
                IF ((fin_giro = '0')) THEN
                    reg_fstate <= Gira_180;
                ELSIF ((fin_giro = '1')) THEN
                    reg_fstate <= Avanza;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Gira_180;
                END IF;

                MD0 <= '0';

                MI0 <= '1';

                MD1 <= '1';

                h_giro <= "10";

                MI1 <= '0';
            WHEN Ganamos =>
                IF ((llego = '0')) THEN
                    reg_fstate <= Avanza;
                ELSIF ((llego = '1')) THEN
                    reg_fstate <= Ganamos;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Ganamos;
                END IF;

                MD0 <= '0';

                MI0 <= '0';

                MD1 <= '0';

                h_giro <= "00";

                MI1 <= '0';
            WHEN OTHERS => 
                MD0 <= 'X';
                MI0 <= 'X';
                MD1 <= 'X';
                MI1 <= 'X';
                h_giro <= "XX";
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
