library verilog;
use verilog.vl_types.all;
entity DFF_fijo_vlg_check_tst is
    port(
        salida          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DFF_fijo_vlg_check_tst;
