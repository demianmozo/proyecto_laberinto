library verilog;
use verilog.vl_types.all;
entity sumador_habilitacion_vlg_vec_tst is
end sumador_habilitacion_vlg_vec_tst;
