-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 07 17:23:46 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LineaRecta IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SR : IN STD_LOGIC := '0';
        SL : IN STD_LOGIC := '0';
        E : IN STD_LOGIC := '0';
        MD0 : OUT STD_LOGIC;
        MI0 : OUT STD_LOGIC;
        MD1 : OUT STD_LOGIC;
        MI1 : OUT STD_LOGIC
    );
END LineaRecta;

ARCHITECTURE BEHAVIOR OF LineaRecta IS
    TYPE type_fstate IS (Idle,Avanza,Dobla_Izquierda,Dobla_Derecha);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= Idle;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,SR,SL,E)
    BEGIN
        MD0 <= '0';
        MI0 <= '0';
        MD1 <= '0';
        MI1 <= '0';
        CASE fstate IS
            WHEN Idle =>
                IF ((E = '1')) THEN
                    reg_fstate <= Avanza;
                ELSIF ((E = '0')) THEN
                    reg_fstate <= Idle;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Idle;
                END IF;

                MD1 <= '0';

                MD0 <= '0';

                MI0 <= '0';

                MI1 <= '0';
            WHEN Avanza =>
                IF ((((E = '1') AND (SR = '0')) AND (SL = '1'))) THEN
                    reg_fstate <= Dobla_Izquierda;
                ELSIF ((((E = '1') AND (SR = '1')) AND (SL = '0'))) THEN
                    reg_fstate <= Dobla_Derecha;
                ELSIF ((((E = '1') AND (SR = '1')) AND (SL = '1'))) THEN
                    reg_fstate <= Avanza;
                ELSIF ((E = '0')) THEN
                    reg_fstate <= Idle;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Avanza;
                END IF;

                MD1 <= '0';

                MD0 <= '1';

                MI0 <= '1';

                MI1 <= '0';
            WHEN Dobla_Izquierda =>
                IF ((((E = '1') AND (SR = '1')) AND (SL = '1'))) THEN
                    reg_fstate <= Avanza;
                ELSIF (((E = '1') AND (SR = '0'))) THEN
                    reg_fstate <= Dobla_Izquierda;
                ELSIF ((E = '0')) THEN
                    reg_fstate <= Idle;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Dobla_Izquierda;
                END IF;

                MD1 <= '0';

                MD0 <= '1';

                MI0 <= '0';

                MI1 <= '1';
            WHEN Dobla_Derecha =>
                IF ((((E = '1') AND (SR = '1')) AND (SL = '1'))) THEN
                    reg_fstate <= Avanza;
                ELSIF (((E = '1') AND (SL = '0'))) THEN
                    reg_fstate <= Dobla_Derecha;
                ELSIF ((E = '0')) THEN
                    reg_fstate <= Idle;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Dobla_Derecha;
                END IF;

                MD1 <= '1';

                MD0 <= '0';

                MI0 <= '1';

                MI1 <= '0';
            WHEN OTHERS => 
                MD0 <= 'X';
                MI0 <= 'X';
                MD1 <= 'X';
                MI1 <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
