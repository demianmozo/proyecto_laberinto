library verilog;
use verilog.vl_types.all;
entity elijo_sentido_vlg_vec_tst is
end elijo_sentido_vlg_vec_tst;
