library verilog;
use verilog.vl_types.all;
entity purbea_vlg_vec_tst is
end purbea_vlg_vec_tst;
