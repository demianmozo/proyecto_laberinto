library verilog;
use verilog.vl_types.all;
entity DFF_fijo_vlg_vec_tst is
end DFF_fijo_vlg_vec_tst;
